module uart(
    input logic        clk,
    input logic        rst,
    input logic        full,

    output logic [7:0] data,
    output logic       wr_en
);



endmodule
